module notgate(
input x,
output y
);
assign y=!x;
endmodule
